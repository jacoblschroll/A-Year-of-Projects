`include "Convolver.v"

// Standard Loop is 10 clock cycles
// 

module A();
    C mod1();
endmodule