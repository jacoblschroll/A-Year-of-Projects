// This handles all operations involving RAM such as read, write, and communication protocols
// Currently this is just a stand in
module memoryController #(parameter addrSize = 14) (clk, rst, address, data);
endmodule